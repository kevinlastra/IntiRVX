

package cpu_configuration;
  parameter xlen = 32;
endpackage
