

package system_config;
  parameter xlen = 64;
endpackage