


package cpu_parameters;

  parameter xlen = 32;
  
endpackage
