

module tb
import pkg::*;
(
  input logic clk,
  input logic rst_n
);

  initial begin
    $display("TEST");
  end

endmodule