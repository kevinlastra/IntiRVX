

package CPU_config;
  parameter xlen = 64;
endpackage