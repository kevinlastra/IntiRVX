
package pkg;

  parameter xlen = 32;
  
endpackage
